module ilevel();

  always @(posedge sum.clk)begin
  $display("block1");
  end
endmodule

module olevel();
  always @(posedge sum.clk)begin
  $display("block2");
  end
endmodule

module top();
     olevel o();
     ilevel i();

endmodule
